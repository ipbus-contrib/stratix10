// (C) 2001-2019 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// -----------------------------------------------
// Reset Synchronizer
// -----------------------------------------------
`timescale 1 ns / 1 ns

module alt_mge_reset_synchronizer
#(
    parameter ASYNC_RESET = 1,
    parameter DEPTH       = 2
)
(
    input   reset_in /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R101" */,

    input   clk,
    output  reset_out
);

    // -----------------------------------------------
    // Synchronizer register chain. We cannot reuse the
    // standard synchronizer in this implementation 
    // because our timing constraints are different.
    //
    // Instead of cutting the timing path to the d-input 
    // on the first flop we need to cut the aclr input.
    // 
    // We omit the "preserve" attribute on the final
    // output register, so that the synthesis tool can
    // duplicate it where needed.
    // -----------------------------------------------
    (*preserve*) reg [DEPTH-1:0] alt_mge_reset_synchronizer_int_chain;
    reg alt_mge_reset_synchronizer_int_chain_out;

    generate if (ASYNC_RESET) begin

        // -----------------------------------------------
        // Assert asynchronously, deassert synchronously.
        // -----------------------------------------------
        always @(posedge clk or posedge reset_in) begin
            if (reset_in) begin
                alt_mge_reset_synchronizer_int_chain <= {DEPTH{1'b1}};
                alt_mge_reset_synchronizer_int_chain_out <= 1'b1;
            end
            else begin
                alt_mge_reset_synchronizer_int_chain[DEPTH-2:0] <= alt_mge_reset_synchronizer_int_chain[DEPTH-1:1];
                alt_mge_reset_synchronizer_int_chain[DEPTH-1] <= 0;
                alt_mge_reset_synchronizer_int_chain_out <= alt_mge_reset_synchronizer_int_chain[0];
            end
        end

        assign reset_out = alt_mge_reset_synchronizer_int_chain_out;
     
    end else begin

        // -----------------------------------------------
        // Assert synchronously, deassert synchronously.
        // -----------------------------------------------
        always @(posedge clk) begin
            alt_mge_reset_synchronizer_int_chain[DEPTH-2:0] <= alt_mge_reset_synchronizer_int_chain[DEPTH-1:1];
            alt_mge_reset_synchronizer_int_chain[DEPTH-1] <= reset_in;
            alt_mge_reset_synchronizer_int_chain_out <= alt_mge_reset_synchronizer_int_chain[0];
        end

        assign reset_out = alt_mge_reset_synchronizer_int_chain_out;
 
    end
    endgenerate

endmodule

