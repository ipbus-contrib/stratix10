package alt_mge_phy_reconfig_parameters_CFG0;

localparam ram_depth = 7;
function [25:0] get_ram_data;
  input integer index;
  automatic reg [0:6][25:0] ram_data = {
    26'h1320400, // [25:16]-DPRIO address=0x132; [15:8]-bit mask=0x04; [2:2]-cdr_pll_set_cdr_vco_speed_fix=60(1'h0);
    26'h1344040, // [25:16]-DPRIO address=0x134; [15:8]-bit mask=0x40; [6:6]-cdr_pll_set_cdr_vco_speed_fix=60(1'h1);
    26'h1354F42, // [25:16]-DPRIO address=0x135; [15:8]-bit mask=0x4F; [6:6]-cdr_pll_set_cdr_vco_speed_fix=60(1'h1); [3:2]-cdr_pll_lf_resistor_pd=lf_pd_setting0(2'h0); [1:0]-cdr_pll_lf_resistor_pfd=lf_pfd_setting2(2'h2);
    26'h1360F0C, // [25:16]-DPRIO address=0x136; [15:8]-bit mask=0x0F; [3:0]-cdr_pll_set_cdr_vco_speed_fix=60(4'hC);
    26'h1390703, // [25:16]-DPRIO address=0x139; [15:8]-bit mask=0x07; [2:0]-cdr_pll_chgpmp_current_pfd=cp_current_pfd_setting3(3'h3);
    26'h13A3F2A, // [25:16]-DPRIO address=0x13A; [15:8]-bit mask=0x3F; [5:3]-cdr_pll_pd_l_counter=8(3'h5); [2:0]-cdr_pll_pfd_l_counter=1(3'h2);
    26'h13BFF28  // [25:16]-DPRIO address=0x13B; [15:8]-bit mask=0xFF; [7:0]-cdr_pll_m_counter=40(8'h28);
};

  begin
  get_ram_data = ram_data[index];
  end
endfunction

localparam PLL_SELECT_VALUE = 1;

localparam HSSI_TX_PLD_PCS_INTERFACE_HD_CHNL_PMA_TX_CLK_HZ_VALUE = 30'd125000000;

localparam HSSI_RX_PLD_PCS_INTERFACE_HD_CHNL_PMA_RX_CLK_HZ_VALUE = 30'd125000000;

localparam PMA_ADAPT_DATARATE_VALUE = "1250000000 bps";

localparam PMA_CGB_DATARATE_VALUE = "1250000000 bps";

localparam PMA_CGB_INPUT_SELECT_X1_VALUE = "lcpll_bot";

localparam PMA_RX_DFE_DATARATE_VALUE = "1250000000 bps";

localparam PMA_RX_ODI_DATARATE_VALUE = "1250000000 bps";

localparam PMA_RX_BUF_DATARATE_VALUE = "1250000000 bps";

localparam PMA_RX_BUF_XRX_PATH_DATARATE_VALUE = "1250000000 bps";

localparam PMA_RX_BUF_XRX_PATH_PMA_RX_DIVCLK_HZ_VALUE = "125000000";

localparam PMA_TX_BUF_DATARATE_VALUE = "1250000000 bps";

localparam PMA_TX_BUF_XTX_PATH_DATARATE_VALUE = "1250000000 bps";

localparam PMA_TX_BUF_XTX_PATH_PMA_TX_DIVCLK_HZ_VALUE = "125000000";

localparam PMA_TX_BUF_XTX_PATH_TX_PLL_CLK_HZ_VALUE = "625000000";

localparam CDR_PLL_DATARATE_VALUE = "1250000000 bps";

localparam CDR_PLL_LPD_COUNTER_VALUE = 5'd8;

localparam CDR_PLL_LPFD_COUNTER_VALUE = 5'd1;

localparam CDR_PLL_OUTPUT_CLOCK_FREQUENCY_VALUE = "625000000 Hz";

localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_VALUE = 8'd60;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_OFST = 306;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD0_OFST = 0;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD0_HIGH = 0;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD0_SIZE = 1;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD0_BITMASK = 32'h00000001;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD0_VALMASK = 32'h00000000;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD0_VALUE = 1'h0;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD1_OFST = 2;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD1_HIGH = 2;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD1_SIZE = 1;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD1_BITMASK = 32'h00000004;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD1_VALMASK = 32'h00000000;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR0_FIELD1_VALUE = 1'h0;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR1_OFST = 308;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR1_FIELD_OFST = 6;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR1_FIELD_HIGH = 6;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR1_FIELD_SIZE = 1;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR1_FIELD_BITMASK = 32'h00000040;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR1_FIELD_VALMASK = 32'h00000040;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR1_FIELD_VALUE = 1'h1;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR2_OFST = 309;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR2_FIELD_OFST = 6;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR2_FIELD_HIGH = 6;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR2_FIELD_SIZE = 1;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR2_FIELD_BITMASK = 32'h00000040;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR2_FIELD_VALMASK = 32'h00000040;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR2_FIELD_VALUE = 1'h1;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR3_OFST = 310;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR3_FIELD_OFST = 0;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR3_FIELD_HIGH = 3;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR3_FIELD_SIZE = 4;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR3_FIELD_BITMASK = 32'h0000000F;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR3_FIELD_VALMASK = 32'h0000000C;
localparam CDR_PLL_SET_CDR_VCO_SPEED_FIX_ADDR3_FIELD_VALUE = 4'hC;

localparam CDR_PLL_VCO_FREQ_VALUE = "5000000000 Hz";

localparam CDR_PLL_CHGPMP_CURRENT_PFD_VALUE = "cp_current_pfd_setting3";
localparam CDR_PLL_CHGPMP_CURRENT_PFD_ADDR_OFST = 313;
localparam CDR_PLL_CHGPMP_CURRENT_PFD_ADDR_FIELD_OFST = 0;
localparam CDR_PLL_CHGPMP_CURRENT_PFD_ADDR_FIELD_HIGH = 2;
localparam CDR_PLL_CHGPMP_CURRENT_PFD_ADDR_FIELD_SIZE = 3;
localparam CDR_PLL_CHGPMP_CURRENT_PFD_ADDR_FIELD_BITMASK = 32'h00000007;
localparam CDR_PLL_CHGPMP_CURRENT_PFD_ADDR_FIELD_VALMASK = 32'h00000003;
localparam CDR_PLL_CHGPMP_CURRENT_PFD_ADDR_FIELD_VALUE = 3'h3;

localparam CDR_PLL_LF_RESISTOR_PD_VALUE = "lf_pd_setting0";
localparam CDR_PLL_LF_RESISTOR_PD_ADDR_OFST = 309;
localparam CDR_PLL_LF_RESISTOR_PD_ADDR_FIELD_OFST = 2;
localparam CDR_PLL_LF_RESISTOR_PD_ADDR_FIELD_HIGH = 3;
localparam CDR_PLL_LF_RESISTOR_PD_ADDR_FIELD_SIZE = 2;
localparam CDR_PLL_LF_RESISTOR_PD_ADDR_FIELD_BITMASK = 32'h0000000C;
localparam CDR_PLL_LF_RESISTOR_PD_ADDR_FIELD_VALMASK = 32'h00000000;
localparam CDR_PLL_LF_RESISTOR_PD_ADDR_FIELD_VALUE = 2'h0;

localparam CDR_PLL_LF_RESISTOR_PFD_VALUE = "lf_pfd_setting2";
localparam CDR_PLL_LF_RESISTOR_PFD_ADDR_OFST = 309;
localparam CDR_PLL_LF_RESISTOR_PFD_ADDR_FIELD_OFST = 0;
localparam CDR_PLL_LF_RESISTOR_PFD_ADDR_FIELD_HIGH = 1;
localparam CDR_PLL_LF_RESISTOR_PFD_ADDR_FIELD_SIZE = 2;
localparam CDR_PLL_LF_RESISTOR_PFD_ADDR_FIELD_BITMASK = 32'h00000003;
localparam CDR_PLL_LF_RESISTOR_PFD_ADDR_FIELD_VALMASK = 32'h00000002;
localparam CDR_PLL_LF_RESISTOR_PFD_ADDR_FIELD_VALUE = 2'h2;

localparam CDR_PLL_M_COUNTER_VALUE = 40;
localparam CDR_PLL_M_COUNTER_ADDR_OFST = 315;
localparam CDR_PLL_M_COUNTER_ADDR_FIELD_OFST = 0;
localparam CDR_PLL_M_COUNTER_ADDR_FIELD_HIGH = 7;
localparam CDR_PLL_M_COUNTER_ADDR_FIELD_SIZE = 8;
localparam CDR_PLL_M_COUNTER_ADDR_FIELD_BITMASK = 32'h000000FF;
localparam CDR_PLL_M_COUNTER_ADDR_FIELD_VALMASK = 32'h00000028;
localparam CDR_PLL_M_COUNTER_ADDR_FIELD_VALUE = 8'h28;

localparam CDR_PLL_PD_L_COUNTER_VALUE = 8;
localparam CDR_PLL_PD_L_COUNTER_ADDR_OFST = 314;
localparam CDR_PLL_PD_L_COUNTER_ADDR_FIELD_OFST = 3;
localparam CDR_PLL_PD_L_COUNTER_ADDR_FIELD_HIGH = 5;
localparam CDR_PLL_PD_L_COUNTER_ADDR_FIELD_SIZE = 3;
localparam CDR_PLL_PD_L_COUNTER_ADDR_FIELD_BITMASK = 32'h00000038;
localparam CDR_PLL_PD_L_COUNTER_ADDR_FIELD_VALMASK = 32'h00000028;
localparam CDR_PLL_PD_L_COUNTER_ADDR_FIELD_VALUE = 3'h5;

localparam CDR_PLL_PFD_L_COUNTER_VALUE = 1;
localparam CDR_PLL_PFD_L_COUNTER_ADDR_OFST = 314;
localparam CDR_PLL_PFD_L_COUNTER_ADDR_FIELD_OFST = 0;
localparam CDR_PLL_PFD_L_COUNTER_ADDR_FIELD_HIGH = 2;
localparam CDR_PLL_PFD_L_COUNTER_ADDR_FIELD_SIZE = 3;
localparam CDR_PLL_PFD_L_COUNTER_ADDR_FIELD_BITMASK = 32'h00000007;
localparam CDR_PLL_PFD_L_COUNTER_ADDR_FIELD_VALMASK = 32'h00000002;
localparam CDR_PLL_PFD_L_COUNTER_ADDR_FIELD_VALUE = 3'h2;

localparam PMA_RX_DESER_DATARATE_VALUE = "1250000000 bps";

endpackage